Stem volume [m3  ha-1] (aboveground) of all trees (in total, per PFT, per Commercial group) on the whole simulated area (average of all hectares).
Time [a1]	Total stem volume [m3 ha-1]	Total Stem Volume per PFT 1 [m3 ha-1]	Total Stem Volume per PFT 2 [m3 ha-1]	Total Stem Volume per PFT 3 [m3 ha-1]	Total Stem Volume per PFT 4 [m3 ha-1]	Total Stem Volume per PFT 5 [m3 ha-1]	Total Stem Volume per PFT 6 [m3 ha-1]	Total stem volume of all non-commercial species [m3 ha-1] 	Total stem volume of all commercial species [m3 ha-1]
Time	TotalStemVolume	StemVolumePerPFT_1	StemVolumePerPFT_2	StemVolumePerPFT_3	StemVolumePerPFT_4	StemVolumePerPFT_5	StemVolumePerPFT_6	StemVolumePerNonCom	StemVolumePerCom
0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00
1.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00	0.000000e+00
2.000000e+00	1.170175e+00	3.701802e-02	2.340449e-01	4.364707e-02	4.232243e-01	3.239877e-03	4.290010e-01	0.000000e+00	1.170175e+00
3.000000e+00	3.006083e+00	7.707779e-02	4.888399e-01	1.192423e-01	9.297555e-01	7.674006e-03	1.383493e+00	0.000000e+00	3.006083e+00
4.000000e+00	6.102254e+00	1.196808e-01	7.902178e-01	2.369199e-01	1.459518e+00	1.362543e-02	3.482293e+00	0.000000e+00	6.102254e+00
5.000000e+00	1.129498e+01	1.707207e-01	1.107440e+00	4.105443e-01	1.899846e+00	1.830368e-02	7.688125e+00	0.000000e+00	1.129498e+01
6.000000e+00	1.997416e+01	2.296913e-01	1.470337e+00	6.791882e-01	2.200312e+00	2.672447e-02	1.536790e+01	0.000000e+00	1.997416e+01
7.000000e+00	3.332706e+01	2.907973e-01	1.861056e+00	1.045980e+00	2.464111e+00	3.586582e-02	2.762925e+01	0.000000e+00	3.332706e+01
8.000000e+00	4.728507e+01	3.465601e-01	2.239786e+00	1.447887e+00	2.714355e+00	4.366004e-02	4.049282e+01	0.000000e+00	4.728507e+01
9.000000e+00	5.910922e+01	4.096963e-01	2.581037e+00	1.930919e+00	2.940838e+00	4.760127e-02	5.119913e+01	0.000000e+00	5.910922e+01
1.000000e+01	6.714088e+01	4.725226e-01	2.959017e+00	2.611168e+00	2.939203e+00	5.418974e-02	5.810478e+01	0.000000e+00	6.714088e+01
1.100000e+01	7.228555e+01	5.361963e-01	3.284080e+00	3.356079e+00	2.913013e+00	6.001476e-02	6.213616e+01	0.000000e+00	7.228555e+01
1.200000e+01	7.803298e+01	6.215784e-01	3.601635e+00	4.394863e+00	2.779221e+00	6.494409e-02	6.657074e+01	0.000000e+00	7.803298e+01
1.300000e+01	8.169498e+01	6.983967e-01	3.877157e+00	5.676775e+00	2.658554e+00	6.295218e-02	6.872114e+01	0.000000e+00	8.169498e+01
1.400000e+01	8.405143e+01	7.873052e-01	4.134996e+00	7.179601e+00	2.578972e+00	6.480180e-02	6.930576e+01	0.000000e+00	8.405143e+01
1.500000e+01	8.558667e+01	8.639176e-01	4.393779e+00	8.986942e+00	2.470241e+00	5.620379e-02	6.881558e+01	0.000000e+00	8.558667e+01
1.600000e+01	8.823481e+01	9.624957e-01	4.687513e+00	1.102316e+01	2.356053e+00	5.992940e-02	6.914566e+01	0.000000e+00	8.823481e+01
1.700000e+01	8.876483e+01	1.060571e+00	4.908013e+00	1.367517e+01	2.246701e+00	4.491572e-02	6.682946e+01	0.000000e+00	8.876483e+01
1.800000e+01	9.003044e+01	1.170911e+00	5.162849e+00	1.607581e+01	2.130818e+00	4.675546e-02	6.544330e+01	0.000000e+00	9.003044e+01
1.900000e+01	9.206898e+01	1.311430e+00	5.501140e+00	1.881450e+01	2.188834e+00	4.862534e-02	6.420445e+01	0.000000e+00	9.206898e+01
2.000000e+01	9.223541e+01	1.437507e+00	5.797384e+00	2.238860e+01	2.223592e+00	5.193789e-02	6.033639e+01	0.000000e+00	9.223541e+01
2.100000e+01	9.192167e+01	1.556068e+00	6.143934e+00	2.501676e+01	2.097069e+00	5.573118e-02	5.705210e+01	0.000000e+00	9.192167e+01
2.200000e+01	9.216633e+01	1.728052e+00	6.553767e+00	2.808400e+01	1.989529e+00	5.842996e-02	5.375256e+01	0.000000e+00	9.216633e+01
2.300000e+01	9.325524e+01	1.902305e+00	6.984594e+00	3.141256e+01	1.894827e+00	6.269166e-02	5.099827e+01	0.000000e+00	9.325524e+01
2.400000e+01	9.307141e+01	2.087679e+00	7.433470e+00	3.401140e+01	2.017057e+00	6.482303e-02	4.745698e+01	0.000000e+00	9.307141e+01
2.500000e+01	9.593110e+01	2.306010e+00	7.951883e+00	3.827276e+01	2.139604e+00	6.853189e-02	4.519231e+01	0.000000e+00	9.593110e+01
2.600000e+01	9.639559e+01	2.550270e+00	8.488678e+00	4.072220e+01	2.027982e+00	6.472505e-02	4.254173e+01	0.000000e+00	9.639559e+01
2.700000e+01	9.949213e+01	2.804710e+00	9.112173e+00	4.477385e+01	1.960983e+00	6.886203e-02	4.077155e+01	0.000000e+00	9.949213e+01
2.800000e+01	1.015615e+02	3.069469e+00	9.817090e+00	4.796947e+01	2.148686e+00	7.468485e-02	3.848214e+01	0.000000e+00	1.015615e+02
2.900000e+01	1.055255e+02	3.360417e+00	1.049638e+01	5.229460e+01	2.055071e+00	7.987848e-02	3.723915e+01	0.000000e+00	1.055255e+02
3.000000e+01	1.087451e+02	3.703792e+00	1.117698e+01	5.630662e+01	1.960608e+00	8.506404e-02	3.551202e+01	0.000000e+00	1.087451e+02
3.100000e+01	1.103551e+02	4.103724e+00	1.188269e+01	5.800818e+01	1.867550e+00	9.227611e-02	3.440063e+01	0.000000e+00	1.103551e+02
3.200000e+01	1.128926e+02	4.504981e+00	1.258797e+01	6.140343e+01	1.778229e+00	9.868001e-02	3.251934e+01	0.000000e+00	1.128926e+02
3.300000e+01	1.167206e+02	4.940271e+00	1.353801e+01	6.486466e+01	1.706105e+00	1.064037e-01	3.156511e+01	0.000000e+00	1.167206e+02
3.400000e+01	1.216422e+02	5.488765e+00	1.452591e+01	6.987555e+01	1.643486e+00	1.137016e-01	2.999475e+01	0.000000e+00	1.216422e+02
3.500000e+01	1.250591e+02	5.940242e+00	1.542035e+01	7.345588e+01	1.549863e+00	1.197682e-01	2.857295e+01	0.000000e+00	1.250591e+02
3.600000e+01	1.269671e+02	6.422841e+00	1.642074e+01	7.593345e+01	1.452036e+00	1.282383e-01	2.660975e+01	0.000000e+00	1.269671e+02
3.700000e+01	1.323661e+02	6.957367e+00	1.715277e+01	8.136385e+01	1.402636e+00	1.372031e-01	2.535230e+01	0.000000e+00	1.323661e+02
3.800000e+01	1.279343e+02	7.586421e+00	1.810763e+01	7.776816e+01	1.304531e+00	1.435369e-01	2.302403e+01	0.000000e+00	1.279343e+02
3.900000e+01	1.323118e+02	8.292196e+00	1.913606e+01	8.157372e+01	1.238039e+00	1.491885e-01	2.192265e+01	0.000000e+00	1.323118e+02
4.000000e+01	1.348058e+02	8.864620e+00	2.027758e+01	8.349437e+01	1.184348e+00	1.576638e-01	2.082727e+01	0.000000e+00	1.348058e+02
4.100000e+01	1.412023e+02	9.712754e+00	2.167562e+01	8.800794e+01	1.129577e+00	1.635231e-01	2.051291e+01	0.000000e+00	1.412023e+02
4.200000e+01	1.435149e+02	1.071483e+01	2.266598e+01	8.916703e+01	1.061581e+00	1.713081e-01	1.973415e+01	0.000000e+00	1.435149e+02
4.300000e+01	1.473031e+02	1.173542e+01	2.392282e+01	9.245798e+01	1.003711e+00	1.785425e-01	1.800458e+01	0.000000e+00	1.473031e+02
4.400000e+01	1.498668e+02	1.258459e+01	2.464412e+01	9.429053e+01	9.502774e-01	1.884349e-01	1.720889e+01	0.000000e+00	1.498668e+02
4.500000e+01	1.565636e+02	1.350659e+01	2.605796e+01	9.915231e+01	9.085475e-01	1.954706e-01	1.674274e+01	0.000000e+00	1.565636e+02
4.600000e+01	1.617706e+02	1.453464e+01	2.723180e+01	1.028155e+02	8.701869e-01	2.010675e-01	1.611744e+01	0.000000e+00	1.617706e+02
4.700000e+01	1.650879e+02	1.550234e+01	2.784325e+01	1.052380e+02	8.138786e-01	2.053793e-01	1.548502e+01	0.000000e+00	1.650879e+02
4.800000e+01	1.701241e+02	1.702067e+01	2.895369e+01	1.083142e+02	7.723579e-01	2.081832e-01	1.485493e+01	0.000000e+00	1.701241e+02
4.900000e+01	1.755260e+02	1.871770e+01	3.022972e+01	1.111025e+02	7.351823e-01	2.081832e-01	1.453277e+01	0.000000e+00	1.755260e+02
5.000000e+01	1.792679e+02	2.031627e+01	3.123607e+01	1.125898e+02	6.995890e-01	2.105346e-01	1.421567e+01	0.000000e+00	1.792679e+02
5.100000e+01	1.763852e+02	2.187889e+01	3.228563e+01	1.078046e+02	6.319412e-01	2.116355e-01	1.357252e+01	0.000000e+00	1.763852e+02
5.200000e+01	1.777710e+02	2.337923e+01	3.397780e+01	1.063541e+02	5.948110e-01	2.128112e-01	1.325228e+01	0.000000e+00	1.777710e+02
5.300000e+01	1.819449e+02	2.569353e+01	3.417584e+01	1.083209e+02	5.705690e-01	2.128112e-01	1.297128e+01	0.000000e+00	1.819449e+02
5.400000e+01	1.875443e+02	2.734244e+01	3.520502e+01	1.118977e+02	5.482422e-01	2.128112e-01	1.233810e+01	0.000000e+00	1.875443e+02
5.500000e+01	1.943997e+02	2.930078e+01	3.620241e+01	1.164461e+02	5.229432e-01	2.128112e-01	1.171467e+01	0.000000e+00	1.943997e+02
5.600000e+01	1.994828e+02	3.183533e+01	3.755687e+01	1.178240e+02	4.979340e-01	2.151626e-01	1.155349e+01	0.000000e+00	1.994828e+02
5.700000e+01	2.045069e+02	3.418832e+01	3.837118e+01	1.198728e+02	4.639035e-01	2.163383e-01	1.139439e+01	0.000000e+00	2.045069e+02
5.800000e+01	2.119654e+02	3.741077e+01	4.055398e+01	1.230307e+02	4.477372e-01	2.151626e-01	1.030705e+01	0.000000e+00	2.119654e+02
5.900000e+01	2.174289e+02	3.942629e+01	4.271908e+01	1.245045e+02	4.191865e-01	2.128112e-01	1.014698e+01	0.000000e+00	2.174289e+02
6.000000e+01	2.272651e+02	4.306010e+01	4.550822e+01	1.285479e+02	4.098872e-01	2.151626e-01	9.523772e+00	0.000000e+00	2.272651e+02
6.100000e+01	2.308940e+02	4.540084e+01	4.699985e+01	1.286824e+02	3.881287e-01	2.151626e-01	9.207575e+00	0.000000e+00	2.308940e+02
6.200000e+01	2.337438e+02	4.738119e+01	4.916218e+01	1.275628e+02	3.696031e-01	2.163383e-01	9.051685e+00	0.000000e+00	2.337438e+02
6.300000e+01	2.399838e+02	5.003925e+01	5.148441e+01	1.294565e+02	3.512821e-01	2.163383e-01	8.435984e+00	0.000000e+00	2.399838e+02
6.400000e+01	2.463113e+02	5.382729e+01	5.274708e+01	1.312193e+02	3.385587e-01	2.151626e-01	7.963901e+00	0.000000e+00	2.463113e+02
6.500000e+01	2.525497e+02	5.826377e+01	5.437669e+01	1.315656e+02	3.206699e-01	2.163383e-01	7.806654e+00	0.000000e+00	2.525497e+02
6.600000e+01	2.478846e+02	6.079093e+01	5.590124e+01	1.233333e+02	3.033498e-01	2.163383e-01	7.339429e+00	0.000000e+00	2.478846e+02
6.700000e+01	2.491368e+02	6.402474e+01	5.839428e+01	1.196526e+02	2.898378e-01	2.175140e-01	6.557876e+00	0.000000e+00	2.491368e+02
6.800000e+01	2.550444e+02	6.921277e+01	5.714815e+01	1.224108e+02	2.744929e-01	2.198654e-01	5.778345e+00	0.000000e+00	2.550444e+02
6.900000e+01	2.645669e+02	7.516200e+01	5.852947e+01	1.250806e+02	2.645797e-01	2.222168e-01	5.308121e+00	0.000000e+00	2.645669e+02
7.000000e+01	2.676478e+02	8.051300e+01	5.958800e+01	1.220734e+02	2.544835e-01	2.233924e-01	4.995499e+00	0.000000e+00	2.676478e+02
7.100000e+01	2.673965e+02	8.042938e+01	5.908190e+01	1.228953e+02	2.377857e-01	2.245681e-01	4.527571e+00	0.000000e+00	2.673965e+02
7.200000e+01	2.634852e+02	8.606274e+01	6.071064e+01	1.118991e+02	2.194685e-01	2.257438e-01	4.367502e+00	0.000000e+00	2.634852e+02
7.300000e+01	2.662095e+02	9.088614e+01	6.107979e+01	1.082514e+02	1.093962e+00	2.233924e-01	4.674781e+00	0.000000e+00	2.662095e+02
7.400000e+01	2.653786e+02	9.249642e+01	6.021305e+01	1.078307e+02	5.385719e-01	2.233924e-01	4.076427e+00	0.000000e+00	2.653786e+02
7.500000e+01	2.711414e+02	9.697880e+01	6.255793e+01	1.067979e+02	5.164485e-01	2.245681e-01	4.065747e+00	0.000000e+00	2.711414e+02
7.600000e+01	2.740071e+02	9.646982e+01	6.451845e+01	1.085495e+02	4.953442e-01	2.269195e-01	3.747104e+00	0.000000e+00	2.740071e+02
7.700000e+01	2.837516e+02	1.027254e+02	6.631587e+01	1.102713e+02	4.745378e-01	2.292709e-01	3.735301e+00	0.000000e+00	2.837516e+02
7.800000e+01	2.871532e+02	1.093441e+02	6.709137e+01	1.064560e+02	4.573407e-01	2.304466e-01	3.573992e+00	0.000000e+00	2.871532e+02
7.900000e+01	2.951348e+02	1.175293e+02	6.948599e+01	1.041928e+02	4.375035e-01	2.304466e-01	3.258798e+00	0.000000e+00	2.951348e+02
8.000000e+01	2.966981e+02	1.196804e+02	7.189743e+01	1.018348e+02	4.200729e-01	2.316223e-01	2.633747e+00	0.000000e+00	2.966981e+02
8.100000e+01	2.929587e+02	1.253112e+02	7.410332e+01	9.060466e+01	4.004107e-01	2.257438e-01	2.313378e+00	0.000000e+00	2.929587e+02
8.200000e+01	2.978317e+02	1.331459e+02	7.314036e+01	8.877959e+01	3.866417e-01	2.280952e-01	2.151099e+00	0.000000e+00	2.978317e+02
8.300000e+01	3.082270e+02	1.403144e+02	7.526920e+01	8.989963e+01	3.691859e-01	2.292709e-01	2.145273e+00	0.000000e+00	3.082270e+02
8.400000e+01	3.196524e+02	1.480955e+02	7.783661e+01	9.101641e+01	3.419510e-01	2.292709e-01	2.132651e+00	0.000000e+00	3.196524e+02
8.500000e+01	3.223514e+02	1.523269e+02	7.835515e+01	8.945116e+01	3.252006e-01	2.257438e-01	1.667249e+00	0.000000e+00	3.223514e+02
8.600000e+01	3.316279e+02	1.623179e+02	7.969851e+01	8.741022e+01	3.129544e-01	2.269195e-01	1.661423e+00	0.000000e+00	3.316279e+02
8.700000e+01	3.300624e+02	1.667752e+02	8.307930e+01	7.817640e+01	3.024571e-01	2.292709e-01	1.499773e+00	0.000000e+00	3.300624e+02
8.800000e+01	3.404393e+02	1.742898e+02	8.532037e+01	7.897753e+01	2.938586e-01	2.250577e-01	1.332650e+00	0.000000e+00	3.404393e+02
8.900000e+01	3.437099e+02	1.818904e+02	8.581979e+01	7.432389e+01	2.801262e-01	2.274091e-01	1.168254e+00	0.000000e+00	3.437099e+02
9.000000e+01	3.546280e+02	1.929378e+02	8.911157e+01	7.091631e+01	2.661770e-01	2.297605e-01	1.166312e+00	0.000000e+00	3.546280e+02
9.100000e+01	3.623692e+02	2.001967e+02	8.898786e+01	7.153612e+01	2.563502e-01	2.297605e-01	1.162428e+00	0.000000e+00	3.623692e+02
9.200000e+01	3.644980e+02	2.094123e+02	8.460120e+01	6.884999e+01	2.450522e-01	2.309362e-01	1.158545e+00	0.000000e+00	3.644980e+02
9.300000e+01	3.722373e+02	2.136312e+02	8.772517e+01	6.940373e+01	2.376820e-01	2.297605e-01	1.009714e+00	0.000000e+00	3.722373e+02
9.400000e+01	3.841951e+02	2.219324e+02	9.082696e+01	6.997246e+01	2.278551e-01	2.285848e-01	1.006801e+00	0.000000e+00	3.841951e+02
9.500000e+01	3.884952e+02	2.303771e+02	9.386313e+01	6.296300e+01	2.155427e-01	2.274091e-01	8.489612e-01	0.000000e+00	3.884952e+02
9.600000e+01	3.952304e+02	2.366563e+02	9.379946e+01	6.349905e+01	2.057158e-01	2.285848e-01	8.411936e-01	0.000000e+00	3.952304e+02
9.700000e+01	4.040124e+02	2.477038e+02	9.527249e+01	5.977780e+01	1.934111e-01	2.285848e-01	8.363389e-01	0.000000e+00	4.040124e+02
9.800000e+01	4.103439e+02	2.547205e+02	9.826385e+01	5.626100e+01	1.884977e-01	2.309362e-01	6.791740e-01	0.000000e+00	4.103439e+02
9.900000e+01	4.071128e+02	2.565162e+02	9.696648e+01	5.254604e+01	1.771837e-01	2.297605e-01	6.772321e-01	0.000000e+00	4.071128e+02
1.000000e+02	4.126005e+02	2.586475e+02	9.994620e+01	5.308447e+01	1.710419e-01	2.297605e-01	5.215707e-01	0.000000e+00	4.126005e+02
1.010000e+02	4.290277e+02	2.715155e+02	1.029795e+02	5.361582e+01	1.661284e-01	2.321119e-01	5.186578e-01	0.000000e+00	4.290277e+02
1.020000e+02	4.271680e+02	2.758044e+02	9.645093e+01	5.415626e+01	1.621702e-01	2.309362e-01	3.633061e-01	0.000000e+00	4.271680e+02
1.030000e+02	4.335493e+02	2.830815e+02	9.369522e+01	5.421301e+01	1.343853e+00	2.368147e-01	9.788849e-01	0.000000e+00	4.335493e+02
1.040000e+02	4.310771e+02	2.850848e+02	9.383370e+01	5.089726e+01	4.905003e-01	2.356390e-01	5.351633e-01	0.000000e+00	4.310771e+02
1.050000e+02	4.473175e+02	2.981926e+02	9.651049e+01	5.137800e+01	4.733032e-01	2.356390e-01	5.273957e-01	0.000000e+00	4.473175e+02
1.060000e+02	4.525285e+02	3.052743e+02	9.421131e+01	5.183648e+01	4.561062e-01	2.344633e-01	5.157444e-01	0.000000e+00	4.525285e+02
1.070000e+02	4.525192e+02	3.079695e+02	9.381957e+01	4.955301e+01	4.401375e-01	2.309362e-01	5.060349e-01	0.000000e+00	4.525192e+02
1.080000e+02	4.331403e+02	2.996493e+02	8.688467e+01	4.545913e+01	4.217121e-01	2.262334e-01	4.992383e-01	0.000000e+00	4.331403e+02
1.090000e+02	4.305678e+02	3.048335e+02	8.232038e+01	4.229214e+01	3.996016e-01	2.297605e-01	4.924417e-01	0.000000e+00	4.305678e+02
1.100000e+02	4.429887e+02	3.146690e+02	8.452752e+01	4.269552e+01	3.873180e-01	2.285848e-01	4.807904e-01	0.000000e+00	4.429887e+02
1.110000e+02	4.549219e+02	3.239900e+02	8.678497e+01	4.306822e+01	3.750344e-01	2.297605e-01	4.739938e-01	0.000000e+00	4.549219e+02
1.120000e+02	4.572850e+02	3.371238e+02	8.004874e+01	3.906029e+01	3.566090e-01	2.274091e-01	4.681681e-01	0.000000e+00	4.572850e+02
1.130000e+02	4.629687e+02	3.439417e+02	7.861100e+01	3.938540e+01	3.406403e-01	2.285848e-01	4.613715e-01	0.000000e+00	4.629687e+02
1.140000e+02	4.720861e+02	3.567103e+02	7.462933e+01	3.974170e+01	3.214736e-01	2.297605e-01	4.536039e-01	0.000000e+00	4.720861e+02
1.150000e+02	4.828277e+02	3.679607e+02	7.561552e+01	3.826576e+01	3.091900e-01	2.297605e-01	4.468073e-01	0.000000e+00	4.828277e+02
1.160000e+02	4.951216e+02	3.810851e+02	7.470434e+01	3.836579e+01	2.956780e-01	2.297605e-01	4.409817e-01	0.000000e+00	4.951216e+02
1.170000e+02	5.006563e+02	3.878495e+02	7.644866e+01	3.540846e+01	2.846228e-01	2.309362e-01	4.341850e-01	0.000000e+00	5.006563e+02
1.180000e+02	5.049087e+02	4.018587e+02	6.914613e+01	3.297426e+01	2.735675e-01	2.285848e-01	4.273884e-01	0.000000e+00	5.049087e+02
1.190000e+02	5.063145e+02	4.021700e+02	7.050045e+01	3.282789e+01	2.023226e-01	2.262334e-01	3.875797e-01	0.000000e+00	5.063145e+02
1.200000e+02	5.095528e+02	4.033040e+02	7.199505e+01	3.308095e+01	4.344828e-01	2.274091e-01	5.108897e-01	0.000000e+00	5.095528e+02
1.210000e+02	5.169212e+02	4.171135e+02	6.529187e+01	3.337028e+01	4.148290e-01	2.285848e-01	5.021512e-01	0.000000e+00	5.169212e+02
1.220000e+02	5.316086e+02	4.313053e+02	6.587096e+01	3.331459e+01	3.988603e-01	2.274091e-01	4.914708e-01	0.000000e+00	5.316086e+02
1.230000e+02	5.406024e+02	4.428974e+02	6.718656e+01	2.943358e+01	3.779782e-01	2.250577e-01	4.817613e-01	0.000000e+00	5.406024e+02
1.240000e+02	5.032588e+02	4.038709e+02	6.851472e+01	2.981401e+01	3.644662e-01	2.227063e-01	4.720519e-01	0.000000e+00	5.032588e+02
1.250000e+02	4.980533e+02	3.969928e+02	6.981246e+01	3.036162e+01	3.534110e-01	2.215307e-01	3.115358e-01	0.000000e+00	4.980533e+02
1.260000e+02	5.092139e+02	4.037745e+02	7.125807e+01	3.079156e+01	1.995729e+00	2.203550e-01	1.173735e+00	0.000000e+00	5.092139e+02
1.270000e+02	5.157967e+02	4.106541e+02	7.254768e+01	3.120291e+01	6.838401e-01	2.180036e-01	4.901896e-01	0.000000e+00	5.157967e+02
1.280000e+02	5.230927e+02	4.213981e+02	7.383502e+01	2.653871e+01	6.371623e-01	2.168279e-01	4.668869e-01	0.000000e+00	5.230927e+02
1.290000e+02	5.373177e+02	4.338204e+02	7.525510e+01	2.696204e+01	6.113668e-01	2.203550e-01	4.484389e-01	0.000000e+00	5.373177e+02
1.300000e+02	5.360607e+02	4.309059e+02	7.652067e+01	2.739259e+01	5.867996e-01	2.180036e-01	4.367876e-01	0.000000e+00	5.360607e+02
1.310000e+02	5.139942e+02	4.110247e+02	7.415036e+01	2.761336e+01	5.671458e-01	2.144765e-01	4.241653e-01	0.000000e+00	5.139942e+02
1.320000e+02	5.054218e+02	3.984772e+02	7.536012e+01	2.808131e+01	2.071888e+00	2.168279e-01	1.214514e+00	0.000000e+00	5.054218e+02
1.330000e+02	5.004660e+02	3.979742e+02	7.630148e+01	2.451805e+01	8.693225e-01	2.156522e-01	5.872840e-01	0.000000e+00	5.004660e+02
1.340000e+02	5.000738e+02	3.992491e+02	7.139552e+01	2.507993e+01	2.652230e+00	2.144765e-01	1.482495e+00	0.000000e+00	5.000738e+02
1.350000e+02	5.046426e+02	4.054219e+02	7.248141e+01	2.468831e+01	1.236560e+00	2.121251e-01	6.022862e-01	0.000000e+00	5.046426e+02
1.360000e+02	5.055324e+02	4.044947e+02	7.377325e+01	2.514226e+01	1.248873e+00	2.121251e-01	6.612231e-01	0.000000e+00	5.055324e+02
1.370000e+02	5.054767e+02	4.114374e+02	6.616869e+01	2.560267e+01	1.266916e+00	2.134652e-01	7.875522e-01	0.000000e+00	5.054767e+02
1.380000e+02	4.939748e+02	3.980357e+02	6.729878e+01	2.609133e+01	1.234347e+00	2.124642e-01	1.102187e+00	0.000000e+00	4.939748e+02
1.390000e+02	5.014760e+02	4.085989e+02	6.309547e+01	2.659733e+01	1.197040e+00	2.138132e-01	1.773411e+00	0.000000e+00	5.014760e+02
1.400000e+02	4.764258e+02	3.816729e+02	6.390879e+01	2.672111e+01	1.067203e+00	2.131549e-01	2.842688e+00	0.000000e+00	4.764258e+02
1.410000e+02	4.892591e+02	3.914290e+02	6.495514e+01	2.732208e+01	9.401047e-01	2.126750e-01	4.400166e+00	0.000000e+00	4.892591e+02
1.420000e+02	4.921789e+02	3.919211e+02	6.608089e+01	2.600383e+01	8.816317e-01	2.147076e-01	7.076788e+00	0.000000e+00	4.921789e+02
1.430000e+02	4.854173e+02	3.854450e+02	6.523238e+01	2.652158e+01	7.711827e-01	2.159154e-01	7.231200e+00	0.000000e+00	4.854173e+02
1.440000e+02	4.899110e+02	3.889485e+02	6.632095e+01	2.705439e+01	9.088627e-01	2.186047e-01	6.459639e+00	0.000000e+00	4.899110e+02
1.450000e+02	4.804265e+02	3.881172e+02	5.875121e+01	2.722023e+01	8.696587e-01	2.217137e-01	5.246470e+00	0.000000e+00	4.804265e+02
1.460000e+02	4.906541e+02	3.974054e+02	5.972630e+01	2.782061e+01	8.368777e-01	2.499957e-01	4.614935e+00	0.000000e+00	4.906541e+02
1.470000e+02	4.872777e+02	3.951581e+02	6.071531e+01	2.621643e+01	7.934263e-01	2.529606e-01	4.141527e+00	0.000000e+00	4.872777e+02
1.480000e+02	4.975028e+02	4.040004e+02	6.184433e+01	2.651029e+01	7.591357e-01	2.567322e-01	4.131817e+00	0.000000e+00	4.975028e+02
1.490000e+02	4.932866e+02	3.989303e+02	6.221681e+01	2.703890e+01	7.193693e-01	2.600071e-01	4.121137e+00	0.000000e+00	4.932866e+02
1.500000e+02	4.923471e+02	4.035347e+02	5.635313e+01	2.753985e+01	6.966964e-01	2.665198e-01	3.956214e+00	0.000000e+00	4.923471e+02
1.510000e+02	4.932030e+02	4.063471e+02	5.665719e+01	2.529948e+01	6.749707e-01	2.739004e-01	3.950388e+00	0.000000e+00	4.932030e+02
1.520000e+02	4.851435e+02	3.941797e+02	5.771432e+01	2.586739e+01	2.397236e+00	2.808500e-01	4.703978e+00	0.000000e+00	4.851435e+02
1.530000e+02	4.923422e+02	4.029222e+02	5.800893e+01	2.650916e+01	9.598684e-01	2.873831e-01	3.654662e+00	0.000000e+00	4.923422e+02
1.540000e+02	4.826243e+02	3.944685e+02	5.889751e+01	2.441021e+01	9.212268e-01	2.945106e-01	3.632330e+00	0.000000e+00	4.826243e+02
1.550000e+02	4.901795e+02	4.004879e+02	5.996552e+01	2.508022e+01	8.847608e-01	3.033753e-01	3.457698e+00	0.000000e+00	4.901795e+02
1.560000e+02	4.600279e+02	3.728436e+02	6.095317e+01	2.194352e+01	8.503667e-01	3.064821e-01	3.130764e+00	0.000000e+00	4.600279e+02
1.570000e+02	4.621553e+02	3.752881e+02	5.989098e+01	2.269819e+01	8.056868e-01	3.171038e-01	3.155246e+00	0.000000e+00	4.621553e+02
1.580000e+02	4.720896e+02	3.832744e+02	6.093738e+01	2.353423e+01	7.756438e-01	3.284583e-01	3.239521e+00	0.000000e+00	4.720896e+02
1.590000e+02	4.817207e+02	3.911358e+02	6.198420e+01	2.403196e+01	7.507953e-01	3.368399e-01	3.481154e+00	0.000000e+00	4.817207e+02
1.600000e+02	4.920940e+02	3.992489e+02	6.299757e+01	2.484314e+01	7.165048e-01	3.444230e-01	3.943498e+00	0.000000e+00	4.920940e+02
1.610000e+02	4.986870e+02	4.038698e+02	6.311257e+01	2.570909e+01	6.618945e-01	3.537923e-01	4.979879e+00	0.000000e+00	4.986870e+02
1.620000e+02	5.037867e+02	4.109701e+02	5.976085e+01	2.568926e+01	5.809263e-01	3.634667e-01	6.422109e+00	0.000000e+00	5.037867e+02
1.630000e+02	5.168263e+02	4.190673e+02	6.074948e+01	2.652703e+01	5.563590e-01	3.729612e-01	9.553204e+00	0.000000e+00	5.168263e+02
1.640000e+02	5.266391e+02	4.270394e+02	6.173256e+01	2.657446e+01	5.293351e-01	3.824481e-01	1.038095e+01	0.000000e+00	5.266391e+02
1.650000e+02	5.275081e+02	4.322816e+02	6.236642e+01	2.260178e+01	5.106285e-01	3.929858e-01	9.354694e+00	0.000000e+00	5.275081e+02
1.660000e+02	5.193266e+02	4.243116e+02	6.336396e+01	2.337889e+01	4.837081e-01	4.009814e-01	7.387452e+00	0.000000e+00	5.193266e+02
1.670000e+02	5.128232e+02	4.133376e+02	6.452210e+01	2.403004e+01	2.631830e+00	2.391661e-01	8.062502e+00	0.000000e+00	5.128232e+02
1.680000e+02	5.106589e+02	4.125090e+02	6.544111e+01	2.486558e+01	8.034667e-01	2.391661e-01	6.800549e+00	0.000000e+00	5.106589e+02
1.690000e+02	5.199771e+02	4.201633e+02	6.655130e+01	2.579207e+01	7.565078e-01	2.393230e-01	6.474587e+00	0.000000e+00	5.199771e+02
1.700000e+02	5.011142e+02	4.118199e+02	5.757447e+01	2.447399e+01	7.080393e-01	2.359683e-01	6.301896e+00	0.000000e+00	5.011142e+02
1.710000e+02	4.959617e+02	4.083509e+02	5.480485e+01	2.363192e+01	2.071520e+00	2.373289e-01	6.865181e+00	0.000000e+00	4.959617e+02
1.720000e+02	5.027182e+02	4.156055e+02	5.528202e+01	2.443630e+01	1.005303e+00	2.364595e-01	6.152645e+00	0.000000e+00	5.027182e+02
1.730000e+02	4.815179e+02	3.947170e+02	5.449634e+01	2.535266e+01	9.153511e-01	2.370359e-01	5.799496e+00	0.000000e+00	4.815179e+02
1.740000e+02	4.906212e+02	4.018172e+02	5.556623e+01	2.633729e+01	8.794474e-01	2.371138e-01	5.783961e+00	0.000000e+00	4.906212e+02
1.750000e+02	4.844751e+02	3.978187e+02	5.571350e+01	2.409377e+01	8.435437e-01	2.372061e-01	5.768426e+00	0.000000e+00	4.844751e+02
1.760000e+02	4.931159e+02	4.048263e+02	5.669246e+01	2.511183e+01	8.046210e-01	2.372557e-01	5.443435e+00	0.000000e+00	4.931159e+02
1.770000e+02	4.808329e+02	3.925048e+02	5.721209e+01	2.484007e+01	7.650322e-01	2.372717e-01	5.273657e+00	0.000000e+00	4.808329e+02
1.780000e+02	4.534098e+02	3.753417e+02	4.885502e+01	2.300311e+01	7.175109e-01	2.372717e-01	5.255209e+00	0.000000e+00	4.534098e+02
1.790000e+02	4.655119e+02	3.817581e+02	4.972992e+01	2.337593e+01	3.828668e+00	2.384829e-01	6.580823e+00	0.000000e+00	4.655119e+02
1.800000e+02	4.646302e+02	3.876508e+02	4.935875e+01	2.122600e+01	1.344641e+00	2.349203e-01	4.815087e+00	0.000000e+00	4.646302e+02
1.810000e+02	4.636415e+02	3.886452e+02	4.814823e+01	2.069265e+01	1.288802e+00	2.349203e-01	4.631716e+00	0.000000e+00	4.636415e+02
1.820000e+02	4.661125e+02	3.896505e+02	4.916107e+01	2.169935e+01	1.235702e+00	7.570145e-02	4.290218e+00	0.000000e+00	4.661125e+02
1.830000e+02	4.638962e+02	3.854486e+02	5.023521e+01	2.284845e+01	1.181372e+00	7.570145e-02	4.106847e+00	0.000000e+00	4.638962e+02
1.840000e+02	4.715832e+02	3.910437e+02	5.133278e+01	2.393426e+01	1.124868e+00	7.570145e-02	4.071893e+00	0.000000e+00	4.715832e+02
1.850000e+02	4.772263e+02	3.975823e+02	4.997426e+01	2.510017e+01	1.069592e+00	7.711407e-02	3.422881e+00	0.000000e+00	4.772263e+02
1.860000e+02	4.567376e+02	3.869979e+02	4.429121e+01	2.110066e+01	1.022914e+00	7.855051e-02	3.246307e+00	0.000000e+00	4.567376e+02
1.870000e+02	4.654159e+02	3.937484e+02	4.528919e+01	2.209055e+01	9.799213e-01	8.002328e-02	3.227859e+00	0.000000e+00	4.654159e+02
1.880000e+02	4.741154e+02	4.000957e+02	4.637840e+01	2.356743e+01	9.430704e-01	8.043144e-02	3.050313e+00	0.000000e+00	4.741154e+02
1.890000e+02	4.796443e+02	4.030787e+02	4.731307e+01	2.523657e+01	9.059384e-01	8.206473e-02	3.027982e+00	0.000000e+00	4.796443e+02
1.900000e+02	4.750785e+02	3.969658e+02	4.836265e+01	2.596666e+01	8.555756e-01	8.130015e-02	2.846552e+00	0.000000e+00	4.750785e+02
1.910000e+02	4.842816e+02	4.034859e+02	4.953625e+01	2.752661e+01	8.196719e-01	8.409910e-02	2.829075e+00	0.000000e+00	4.842816e+02
1.920000e+02	4.838223e+02	4.034274e+02	5.046898e+01	2.659278e+01	7.533405e-01	8.635485e-02	2.493403e+00	0.000000e+00	4.838223e+02
1.930000e+02	4.875208e+02	4.063761e+02	5.081955e+01	2.703245e+01	7.275449e-01	8.532936e-02	2.479810e+00	0.000000e+00	4.875208e+02
1.940000e+02	4.775024e+02	4.128959e+02	4.121780e+01	2.016672e+01	6.793576e-01	8.702852e-02	2.455537e+00	0.000000e+00	4.775024e+02
1.950000e+02	4.682030e+02	4.014368e+02	4.201147e+01	2.172344e+01	6.535620e-01	8.904217e-02	2.288672e+00	0.000000e+00	4.682030e+02
1.960000e+02	4.690420e+02	3.999449e+02	4.303683e+01	2.322570e+01	6.213435e-01	9.046670e-02	2.122778e+00	0.000000e+00	4.690420e+02
1.970000e+02	4.598600e+02	3.909991e+02	4.311789e+01	2.310130e+01	5.903532e-01	9.351509e-02	1.957854e+00	0.000000e+00	4.598600e+02
1.980000e+02	4.681354e+02	3.972490e+02	4.418578e+01	2.424234e+01	5.667332e-01	9.951713e-02	1.791960e+00	0.000000e+00	4.681354e+02
1.990000e+02	4.770201e+02	4.035798e+02	4.550298e+01	2.566408e+01	5.384809e-01	1.038123e-01	1.630921e+00	0.000000e+00	4.770201e+02
2.000000e+02	4.719508e+02	3.990153e+02	4.381657e+01	2.704612e+01	5.040868e-01	1.085189e-01	1.460172e+00	0.000000e+00	4.719508e+02
2.010000e+02	4.817772e+02	4.049933e+02	4.455716e+01	2.623315e+01	3.192969e+00	8.290146e-02	2.717683e+00	0.000000e+00	4.817772e+02
2.020000e+02	4.815744e+02	4.103267e+02	4.088407e+01	2.798814e+01	8.210039e-01	8.055007e-02	1.473903e+00	0.000000e+00	4.815744e+02
2.030000e+02	4.899333e+02	4.164874e+02	4.190175e+01	2.922082e+01	7.853814e-01	8.055007e-02	1.457397e+00	0.000000e+00	4.899333e+02
2.040000e+02	4.971500e+02	4.233706e+02	4.107128e+01	3.058893e+01	7.531628e-01	7.937438e-02	1.286648e+00	0.000000e+00	4.971500e+02
2.050000e+02	5.060519e+02	4.292010e+02	4.221704e+01	3.286864e+01	7.249105e-01	8.055007e-02	9.597144e-01	0.000000e+00	5.060519e+02
2.060000e+02	5.079493e+02	4.291731e+02	4.331662e+01	3.374513e+01	6.914636e-01	8.172577e-02	9.412665e-01	0.000000e+00	5.079493e+02
2.070000e+02	4.713870e+02	3.942942e+02	4.114326e+01	3.432057e+01	6.423291e-01	7.937438e-02	9.072834e-01	0.000000e+00	4.713870e+02
2.080000e+02	4.841394e+02	4.012845e+02	4.130050e+01	3.587639e+01	3.401228e+00	7.702299e-02	2.199748e+00	0.000000e+00	4.841394e+02
2.090000e+02	4.870848e+02	4.054856e+02	4.212630e+01	3.751545e+01	9.629313e-01	7.349591e-02	9.210141e-01	0.000000e+00	4.870848e+02
2.100000e+02	4.926227e+02	4.088280e+02	4.299964e+01	3.890398e+01	9.144628e-01	7.702299e-02	8.996533e-01	0.000000e+00	4.926227e+02
2.110000e+02	5.007812e+02	4.147338e+02	4.384521e+01	4.036893e+01	8.763837e-01	7.467160e-02	8.821763e-01	0.000000e+00	5.007812e+02
2.120000e+02	4.696535e+02	3.873930e+02	4.094805e+01	3.953278e+01	8.444463e-01	7.349591e-02	8.617865e-01	0.000000e+00	4.696535e+02
2.130000e+02	4.758501e+02	3.868484e+02	4.185628e+01	4.113179e+01	3.620542e+00	7.584730e-02	2.317232e+00	0.000000e+00	4.758501e+02
2.140000e+02	4.734119e+02	3.866597e+02	4.227261e+01	4.224984e+01	1.140481e+00	7.702299e-02	1.012283e+00	0.000000e+00	4.734119e+02
2.150000e+02	4.633423e+02	3.784950e+02	4.314803e+01	3.954993e+01	1.086433e+00	8.172577e-02	9.812126e-01	0.000000e+00	4.633423e+02
2.160000e+02	4.702719e+02	3.849724e+02	4.369241e+01	3.953513e+01	1.032385e+00	8.172577e-02	9.579100e-01	0.000000e+00	4.702719e+02
2.170000e+02	4.795142e+02	3.912000e+02	4.464293e+01	4.166044e+01	9.906212e-01	8.172577e-02	9.384911e-01	0.000000e+00	4.795142e+02
2.180000e+02	4.878484e+02	3.965932e+02	4.555748e+01	4.390756e+01	9.451719e-01	8.407716e-02	7.609457e-01	0.000000e+00	4.878484e+02
2.190000e+02	4.930592e+02	4.035864e+02	4.623054e+01	4.154558e+01	8.825255e-01	8.525285e-02	7.289045e-01	0.000000e+00	4.930592e+02
2.200000e+02	4.949604e+02	4.075243e+02	4.399739e+01	4.180803e+01	8.395328e-01	8.362018e-02	7.075437e-01	0.000000e+00	4.949604e+02
2.210000e+02	4.626917e+02	3.890328e+02	3.694072e+01	3.513181e+01	8.088238e-01	8.362018e-02	6.939505e-01	0.000000e+00	4.626917e+02
2.220000e+02	4.666723e+02	3.930538e+02	3.772376e+01	3.435895e+01	7.756581e-01	8.362018e-02	6.764735e-01	0.000000e+00	4.666723e+02
2.230000e+02	4.726769e+02	3.979550e+02	3.879521e+01	3.443228e+01	7.486341e-01	8.479588e-02	6.609384e-01	0.000000e+00	4.726769e+02
2.240000e+02	4.764352e+02	4.032030e+02	3.934414e+01	3.244919e+01	7.154684e-01	8.479588e-02	6.386066e-01	0.000000e+00	4.764352e+02
2.250000e+02	4.847330e+02	4.106273e+02	3.967377e+01	3.304346e+01	6.847594e-01	8.362018e-02	6.201587e-01	0.000000e+00	4.847330e+02
2.260000e+02	4.605348e+02	3.836443e+02	4.090764e+01	3.478660e+01	6.601922e-01	8.479588e-02	4.513518e-01	0.000000e+00	4.605348e+02
2.270000e+02	4.722813e+02	3.912784e+02	3.876901e+01	3.642126e+01	3.688102e+00	8.479588e-02	2.039817e+00	0.000000e+00	4.722813e+02
2.280000e+02	4.764919e+02	3.967934e+02	3.974932e+01	3.650349e+01	2.139139e+00	8.126879e-02	1.225195e+00	0.000000e+00	4.764919e+02
2.290000e+02	4.846091e+02	4.045068e+02	3.983946e+01	3.818223e+01	1.246120e+00	8.027739e-02	7.542865e-01	0.000000e+00	4.846091e+02
2.300000e+02	4.920968e+02	4.120168e+02	3.992228e+01	3.815363e+01	1.195476e+00	8.048006e-02	7.280710e-01	0.000000e+00	4.920968e+02
2.310000e+02	4.788561e+02	3.975989e+02	4.076660e+01	3.872863e+01	1.141428e+00	8.068679e-02	5.398452e-01	0.000000e+00	4.788561e+02
2.320000e+02	4.794748e+02	3.968108e+02	4.049779e+01	4.046773e+01	1.095979e+00	8.207335e-02	5.204263e-01	0.000000e+00	4.794748e+02
2.330000e+02	4.886633e+02	4.050489e+02	4.085723e+01	4.112454e+01	1.051758e+00	8.466574e-02	4.961527e-01	0.000000e+00	4.886633e+02
2.340000e+02	4.677035e+02	3.858232e+02	4.151196e+01	3.883290e+01	9.866549e-01	8.378472e-02	4.650824e-01	0.000000e+00	4.677035e+02
2.350000e+02	4.823675e+02	3.943067e+02	4.213118e+01	3.957756e+01	4.143542e+00	8.408684e-02	2.124427e+00	0.000000e+00	4.823675e+02
2.360000e+02	4.633898e+02	3.784059e+02	4.199003e+01	4.098884e+01	1.310572e+00	7.986146e-02	6.146079e-01	0.000000e+00	4.633898e+02
2.370000e+02	4.718236e+02	3.816922e+02	4.302966e+01	4.012383e+01	4.545431e+00	8.184970e-02	2.350636e+00	0.000000e+00	4.718236e+02
2.380000e+02	4.638081e+02	3.776364e+02	4.341518e+01	4.014405e+01	1.707716e+00	5.702341e-02	8.478080e-01	0.000000e+00	4.638081e+02
2.390000e+02	4.654794e+02	3.844942e+02	4.311085e+01	3.519253e+01	1.678230e+00	5.998452e-02	9.436117e-01	0.000000e+00	4.654794e+02
2.400000e+02	4.755744e+02	3.924201e+02	4.365153e+01	3.655682e+01	1.647877e+00	6.181501e-02	1.236278e+00	0.000000e+00	4.755744e+02
2.410000e+02	4.877220e+02	4.016347e+02	4.471311e+01	3.787985e+01	1.575236e+00	6.124660e-02	1.857903e+00	0.000000e+00	4.877220e+02
2.420000e+02	4.544478e+02	3.842843e+02	2.695205e+01	3.885463e+01	1.429145e+00	6.151270e-02	2.866221e+00	0.000000e+00	4.544478e+02
2.430000e+02	4.745091e+02	3.929171e+02	2.809721e+01	3.516951e+01	9.574258e+00	6.180011e-02	8.689202e+00	0.000000e+00	4.745091e+02
2.440000e+02	4.396840e+02	3.661961e+02	2.886384e+01	3.443628e+01	2.297526e+00	6.145362e-02	7.828719e+00	0.000000e+00	4.396840e+02
2.450000e+02	4.163745e+02	3.461727e+02	2.434148e+01	3.602789e+01	2.181218e+00	6.629358e-02	7.584847e+00	0.000000e+00	4.163745e+02
2.460000e+02	4.269434e+02	3.549793e+02	2.548749e+01	3.728481e+01	2.086942e+00	7.374859e-02	7.031107e+00	0.000000e+00	4.269434e+02
2.470000e+02	4.104914e+02	3.420919e+02	2.575261e+01	3.493119e+01	1.987752e+00	7.767312e-02	5.650277e+00	0.000000e+00	4.104914e+02
2.480000e+02	4.015666e+02	3.322263e+02	2.692764e+01	3.513807e+01	1.898160e+00	7.959935e-02	5.296862e+00	0.000000e+00	4.015666e+02
2.490000e+02	4.120249e+02	3.422426e+02	2.656468e+01	3.672319e+01	1.795285e+00	7.996552e-02	4.619160e+00	0.000000e+00	4.120249e+02
2.500000e+02	4.061228e+02	3.416326e+02	2.626448e+01	3.185092e+01	1.708917e+00	8.167096e-02	4.584206e+00	0.000000e+00	4.061228e+02
2.510000e+02	4.138672e+02	3.519003e+02	2.743999e+01	2.860225e+01	1.614489e+00	7.260219e-02	4.237587e+00	0.000000e+00	4.138672e+02
2.520000e+02	4.179780e+02	3.555562e+02	2.707167e+01	3.018724e+01	1.510003e+00	7.260219e-02	3.580275e+00	0.000000e+00	4.179780e+02
2.530000e+02	4.308628e+02	3.661669e+02	2.778992e+01	3.184592e+01	1.439834e+00	7.495358e-02	3.545321e+00	0.000000e+00	4.308628e+02
2.540000e+02	4.432910e+02	3.759803e+02	2.897966e+01	3.335873e+01	1.382869e+00	7.612928e-02	3.513280e+00	0.000000e+00	4.432910e+02
2.550000e+02	4.487895e+02	3.818590e+02	2.830757e+01	3.404627e+01	1.327133e+00	7.612928e-02	3.173458e+00	0.000000e+00	4.487895e+02
2.560000e+02	4.624653e+02	3.929913e+02	2.941911e+01	3.572745e+01	1.266713e+00	7.612928e-02	2.984614e+00	0.000000e+00	4.624653e+02
2.570000e+02	4.627264e+02	3.912613e+02	3.047169e+01	3.697084e+01	1.167984e+00	7.730497e-02	2.777322e+00	0.000000e+00	4.627264e+02
2.580000e+02	4.707337e+02	4.008911e+02	3.072312e+01	3.516036e+01	1.128676e+00	7.730497e-02	2.753048e+00	0.000000e+00	4.707337e+02
2.590000e+02	4.810549e+02	4.122255e+02	2.845454e+01	3.696722e+01	1.066415e+00	7.320719e-02	2.268074e+00	0.000000e+00	4.810549e+02
2.600000e+02	4.914564e+02	4.230181e+02	2.959803e+01	3.549039e+01	1.021964e+00	7.438288e-02	2.253510e+00	0.000000e+00	4.914564e+02
2.610000e+02	5.007045e+02	4.312489e+02	2.885892e+01	3.731993e+01	9.760544e-01	7.438288e-02	2.226324e+00	0.000000e+00	5.007045e+02
2.620000e+02	5.129292e+02	4.433155e+02	2.993472e+01	3.646134e+01	9.414301e-01	7.320719e-02	2.203021e+00	0.000000e+00	5.129292e+02
2.630000e+02	5.139923e+02	4.431852e+02	3.032399e+01	3.710649e+01	1.245833e+00	6.850441e-02	2.062243e+00	0.000000e+00	5.139923e+02
2.640000e+02	5.163595e+02	4.463495e+02	3.118344e+01	3.565596e+01	1.098048e+00	7.438288e-02	1.998160e+00	0.000000e+00	5.163595e+02
2.650000e+02	5.050737e+02	4.325532e+02	3.203652e+01	3.738065e+01	1.052368e+00	7.320719e-02	1.977770e+00	0.000000e+00	5.050737e+02
2.660000e+02	5.096758e+02	4.339391e+02	3.163034e+01	3.569470e+01	4.633808e+00	7.320719e-02	3.704600e+00	0.000000e+00	5.096758e+02
2.670000e+02	5.123505e+02	4.400476e+02	3.222442e+01	3.667752e+01	1.349077e+00	7.555858e-02	1.976318e+00	0.000000e+00	5.123505e+02
2.680000e+02	5.158450e+02	4.407354e+02	3.337993e+01	3.846447e+01	1.329453e+00	7.673427e-02	1.859023e+00	0.000000e+00	5.158450e+02
2.690000e+02	5.289343e+02	4.515433e+02	3.393739e+01	4.013800e+01	1.366637e+00	7.673427e-02	1.872159e+00	0.000000e+00	5.289343e+02
2.700000e+02	5.263016e+02	4.542794e+02	3.099512e+01	3.758283e+01	1.366212e+00	7.790997e-02	2.000106e+00	0.000000e+00	5.263016e+02
2.710000e+02	5.411008e+02	4.662548e+02	3.177535e+01	3.928035e+01	1.367632e+00	7.790997e-02	2.344779e+00	0.000000e+00	5.411008e+02
2.720000e+02	5.461164e+02	4.681406e+02	3.261745e+01	4.091774e+01	1.333399e+00	7.673427e-02	3.030500e+00	0.000000e+00	5.461164e+02
2.730000e+02	5.366859e+02	4.582964e+02	3.337475e+01	3.977227e+01	1.166181e+00	7.438288e-02	4.001948e+00	0.000000e+00	5.366859e+02
2.740000e+02	5.422512e+02	4.625174e+02	3.439653e+01	3.913868e+01	1.030980e+00	7.438288e-02	5.093281e+00	0.000000e+00	5.422512e+02
2.750000e+02	5.522893e+02	4.722851e+02	3.512577e+01	3.658079e+01	9.394982e-01	7.555858e-02	7.282577e+00	0.000000e+00	5.522893e+02
2.760000e+02	5.678918e+02	4.843192e+02	3.618590e+01	3.795812e+01	8.933682e-01	7.085580e-02	8.464368e+00	0.000000e+00	5.678918e+02
2.770000e+02	5.730952e+02	4.920860e+02	3.553465e+01	3.705154e+01	8.519216e-01	7.085580e-02	7.500256e+00	0.000000e+00	5.730952e+02
2.780000e+02	5.756774e+02	4.943155e+02	3.581889e+01	3.836732e+01	8.328687e-01	7.320719e-02	6.269682e+00	0.000000e+00	5.756774e+02
2.790000e+02	5.691281e+02	4.886925e+02	3.668835e+01	3.692679e+01	7.971665e-01	7.438288e-02	5.948927e+00	0.000000e+00	5.691281e+02
2.800000e+02	5.707606e+02	4.931867e+02	3.462020e+01	3.651656e+01	7.356953e-01	7.555858e-02	5.625877e+00	0.000000e+00	5.707606e+02
2.810000e+02	5.688738e+02	4.888328e+02	3.580092e+01	3.783644e+01	7.077872e-01	7.673427e-02	5.619081e+00	0.000000e+00	5.688738e+02
2.820000e+02	5.698269e+02	4.891761e+02	3.690935e+01	3.768443e+01	6.844484e-01	7.555858e-02	5.297002e+00	0.000000e+00	5.698269e+02
2.830000e+02	5.677319e+02	4.851238e+02	3.810631e+01	3.879737e+01	6.456886e-01	8.378844e-02	4.974923e+00	0.000000e+00	5.677319e+02
2.840000e+02	5.771785e+02	4.940108e+02	3.761863e+01	4.002721e+01	6.241524e-01	8.378844e-02	4.813884e+00	0.000000e+00	5.771785e+02
2.850000e+02	5.862374e+02	5.012821e+02	3.813247e+01	4.133236e+01	5.995586e-01	8.378844e-02	4.807087e+00	0.000000e+00	5.862374e+02
2.860000e+02	5.799565e+02	4.950743e+02	3.724868e+01	4.216731e+01	5.811332e-01	8.378844e-02	4.801262e+00	0.000000e+00	5.799565e+02
2.870000e+02	5.558776e+02	4.752568e+02	3.787171e+01	3.750112e+01	5.332006e-01	8.231423e-02	4.632455e+00	0.000000e+00	5.558776e+02
2.880000e+02	5.616308e+02	4.782658e+02	3.914190e+01	3.832285e+01	1.157809e+00	8.701701e-02	4.655414e+00	0.000000e+00	5.616308e+02
2.890000e+02	5.609232e+02	4.764667e+02	3.989915e+01	3.947631e+01	8.212379e-01	9.054409e-02	4.169245e+00	0.000000e+00	5.609232e+02
2.900000e+02	5.480479e+02	4.615728e+02	4.056026e+01	4.089166e+01	7.757354e-01	9.171979e-02	4.155652e+00	0.000000e+00	5.480479e+02
2.910000e+02	5.597349e+02	4.716611e+02	4.105086e+01	4.235111e+01	7.443724e-01	9.289548e-02	3.834544e+00	0.000000e+00	5.597349e+02
2.920000e+02	5.714859e+02	4.819154e+02	4.225533e+01	4.300732e+01	7.084932e-01	9.171979e-02	3.507611e+00	0.000000e+00	5.714859e+02
2.930000e+02	5.505861e+02	4.642059e+02	4.173089e+01	4.089587e+01	6.476495e-01	8.936840e-02	3.016459e+00	0.000000e+00	5.505861e+02
2.940000e+02	5.459339e+02	4.587309e+02	4.249863e+01	4.133670e+01	5.935219e-01	9.054409e-02	2.683700e+00	0.000000e+00	5.459339e+02
2.950000e+02	5.517661e+02	4.683963e+02	4.067306e+01	3.952293e+01	5.615579e-01	9.054409e-02	2.521690e+00	0.000000e+00	5.517661e+02
2.960000e+02	5.512232e+02	4.709465e+02	3.846861e+01	3.865644e+01	5.429024e-01	9.289548e-02	2.515864e+00	0.000000e+00	5.512232e+02
2.970000e+02	5.612856e+02	4.807315e+02	3.809011e+01	3.934804e+01	5.195369e-01	8.936840e-02	2.507125e+00	0.000000e+00	5.612856e+02
2.980000e+02	5.591799e+02	4.814749e+02	3.903816e+01	3.589519e+01	4.949432e-01	8.936840e-02	2.187341e+00	0.000000e+00	5.591799e+02
2.990000e+02	5.664328e+02	4.903101e+02	4.008857e+01	3.328272e+01	4.789745e-01	9.289548e-02	2.179573e+00	0.000000e+00	5.664328e+02
3.000000e+02	5.658985e+02	4.878302e+02	4.119705e+01	3.414105e+01	4.633765e-01	9.407118e-02	2.172777e+00	0.000000e+00	5.658985e+02
3.010000e+02	5.531833e+02	4.732911e+02	4.200118e+01	3.518298e+01	4.486362e-01	9.642257e-02	2.163067e+00	0.000000e+00	5.531833e+02
3.020000e+02	5.191025e+02	4.415119e+02	3.863004e+01	3.627364e+01	4.357251e-01	9.877396e-02	2.152387e+00	0.000000e+00	5.191025e+02
3.030000e+02	5.304452e+02	4.506318e+02	3.970042e+01	3.745200e+01	4.148164e-01	9.759826e-02	2.148503e+00	0.000000e+00	5.304452e+02
3.040000e+02	5.272810e+02	4.475450e+02	4.063941e+01	3.670470e+01	3.404873e-01	9.407118e-02	1.957365e+00	0.000000e+00	5.272810e+02
3.050000e+02	5.289623e+02	4.566651e+02	3.479018e+01	3.492910e+01	5.603373e-01	9.407118e-02	1.923519e+00	0.000000e+00	5.289623e+02
3.060000e+02	5.296253e+02	4.559362e+02	3.552420e+01	3.577278e+01	5.382003e-01	9.407118e-02	1.759919e+00	0.000000e+00	5.296253e+02
3.070000e+02	5.383400e+02	4.648832e+02	3.570774e+01	3.539350e+01	5.136065e-01	9.171979e-02	1.750210e+00	0.000000e+00	5.383400e+02
3.080000e+02	5.129985e+02	4.382955e+02	3.623055e+01	3.630570e+01	4.933252e-01	8.819270e-02	1.585287e+00	0.000000e+00	5.129985e+02
3.090000e+02	5.257425e+02	4.462764e+02	3.709023e+01	3.726063e+01	2.426138e+00	8.819270e-02	2.600895e+00	0.000000e+00	5.257425e+02
3.100000e+02	5.098442e+02	4.311966e+02	3.791253e+01	3.807478e+01	8.126725e-01	8.466562e-02	1.762969e+00	0.000000e+00	5.098442e+02
3.110000e+02	5.100289e+02	4.396516e+02	3.515284e+01	3.277699e+01	7.776509e-01	8.348992e-02	1.586395e+00	0.000000e+00	5.100289e+02
3.120000e+02	5.112206e+02	4.473754e+02	3.150226e+01	2.993744e+01	7.491685e-01	8.348992e-02	1.572802e+00	0.000000e+00	5.112206e+02
3.130000e+02	5.003082e+02	4.363505e+02	3.099025e+01	3.070276e+01	6.478154e-01	8.584131e-02	1.531051e+00	0.000000e+00	5.003082e+02
3.140000e+02	5.046865e+02	4.424634e+02	3.074880e+01	2.939879e+01	6.257049e-01	8.466562e-02	1.365157e+00	0.000000e+00	5.046865e+02
3.150000e+02	5.100856e+02	4.486839e+02	3.150384e+01	2.785561e+01	6.017386e-01	8.701701e-02	1.353506e+00	0.000000e+00	5.100856e+02
3.160000e+02	5.133026e+02	4.517987e+02	3.194780e+01	2.785290e+01	5.814574e-01	8.936840e-02	1.032398e+00	0.000000e+00	5.133026e+02
3.170000e+02	4.732639e+02	4.192247e+02	2.707665e+01	2.530998e+01	5.507483e-01	8.008058e-02	1.021717e+00	0.000000e+00	4.732639e+02
3.180000e+02	4.687336e+02	4.160113e+02	2.325527e+01	2.609773e+01	1.683297e+00	7.786042e-02	1.608168e+00	0.000000e+00	4.687336e+02
3.190000e+02	4.834517e+02	4.238644e+02	2.387598e+01	2.690749e+01	5.251685e+00	7.290867e-02	3.479178e+00	0.000000e+00	4.834517e+02
3.200000e+02	4.849959e+02	4.303072e+02	2.434802e+01	2.768952e+01	1.215292e+00	7.437855e-02	1.361548e+00	0.000000e+00	4.849959e+02
3.210000e+02	4.867341e+02	4.334125e+02	2.495715e+01	2.578864e+01	1.163700e+00	7.584103e-02	1.336303e+00	0.000000e+00	4.867341e+02
3.220000e+02	4.734295e+02	4.220293e+02	2.233763e+01	2.655706e+01	1.117624e+00	7.877112e-02	1.309117e+00	0.000000e+00	4.734295e+02
3.230000e+02	4.858822e+02	4.293978e+02	2.299282e+01	2.697864e+01	3.747544e+00	8.043849e-02	2.684945e+00	0.000000e+00	4.858822e+02
3.240000e+02	4.914816e+02	4.373153e+02	2.351355e+01	2.772373e+01	1.394376e+00	8.089867e-02	1.453788e+00	0.000000e+00	4.914816e+02
3.250000e+02	4.848463e+02	4.294195e+02	2.417689e+01	2.855554e+01	1.340328e+00	8.366825e-02	1.270417e+00	0.000000e+00	4.848463e+02
3.260000e+02	4.984491e+02	4.354724e+02	2.431899e+01	2.925327e+01	5.744001e+00	8.398258e-02	3.576410e+00	0.000000e+00	4.984491e+02
3.270000e+02	4.878904e+02	4.333144e+02	2.462053e+01	2.686096e+01	1.606882e+00	8.222172e-02	1.405378e+00	0.000000e+00	4.878904e+02
3.280000e+02	4.905046e+02	4.407540e+02	2.002261e+01	2.690125e+01	1.536238e+00	7.815184e-02	1.212297e+00	0.000000e+00	4.905046e+02
3.290000e+02	4.898884e+02	4.392305e+02	2.050178e+01	2.743000e+01	1.469906e+00	7.880059e-02	1.177343e+00	0.000000e+00	4.898884e+02
3.300000e+02	4.940489e+02	4.467215e+02	1.784840e+01	2.700755e+01	1.401719e+00	7.959759e-02	9.900886e-01	0.000000e+00	4.940489e+02
3.310000e+02	5.028445e+02	4.542932e+02	1.818725e+01	2.797362e+01	1.346443e+00	8.306194e-02	9.609602e-01	0.000000e+00	5.028445e+02
3.320000e+02	4.945845e+02	4.454176e+02	1.869168e+01	2.835966e+01	1.149278e+00	7.607529e-02	8.901822e-01	0.000000e+00	4.945845e+02
3.330000e+02	4.897645e+02	4.391548e+02	1.909934e+01	2.926001e+01	1.204554e+00	7.489960e-02	9.708723e-01	0.000000e+00	4.897645e+02
3.340000e+02	4.752890e+02	4.230889e+02	1.958559e+01	3.031808e+01	1.154191e+00	7.287098e-02	1.069397e+00	0.000000e+00	4.752890e+02
3.350000e+02	4.869039e+02	4.305731e+02	2.022121e+01	3.094339e+01	2.833360e+00	7.440619e-02	2.258443e+00	0.000000e+00	4.869039e+02
3.360000e+02	4.824484e+02	4.265496e+02	2.051207e+01	3.211067e+01	1.382666e+00	7.463178e-02	1.818742e+00	0.000000e+00	4.824484e+02
3.370000e+02	4.918482e+02	4.338812e+02	2.119435e+01	3.263199e+01	1.328618e+00	7.580747e-02	2.736200e+00	0.000000e+00	4.918482e+02
3.380000e+02	5.001289e+02	4.412521e+02	1.934959e+01	3.381913e+01	1.263515e+00	7.463178e-02	4.369998e+00	0.000000e+00	5.001289e+02
3.390000e+02	5.088057e+02	4.458479e+02	1.990672e+01	3.517091e+01	1.198386e+00	7.815886e-02	6.603625e+00	0.000000e+00	5.088057e+02
3.400000e+02	5.178132e+02	4.532513e+02	2.056135e+01	3.580517e+01	1.146794e+00	7.933455e-02	6.969205e+00	0.000000e+00	5.178132e+02
3.410000e+02	5.228834e+02	4.607078e+02	2.121053e+01	3.380659e+01	1.094576e+00	7.815886e-02	5.985770e+00	0.000000e+00	5.228834e+02
3.420000e+02	5.224098e+02	4.605240e+02	2.162193e+01	3.443792e+01	1.054040e+00	7.815886e-02	4.693751e+00	0.000000e+00	5.224098e+02
3.430000e+02	5.310914e+02	4.679819e+02	2.158222e+01	3.608344e+01	9.993645e-01	7.815886e-02	4.366319e+00	0.000000e+00	5.310914e+02
3.440000e+02	5.242583e+02	4.596734e+02	2.163550e+01	3.789596e+01	9.446892e-01	7.815886e-02	4.030587e+00	0.000000e+00	5.242583e+02
3.450000e+02	5.274338e+02	4.622509e+02	2.221222e+01	3.797931e+01	9.016965e-01	7.657916e-02	4.013110e+00	0.000000e+00	5.274338e+02
3.460000e+02	4.931130e+02	4.319555e+02	2.097197e+01	3.549642e+01	8.009710e-01	7.422777e-02	3.813862e+00	0.000000e+00	4.931130e+02
3.470000e+02	4.935543e+02	4.254389e+02	2.139353e+01	3.427508e+01	5.988940e+00	7.540347e-02	6.382431e+00	0.000000e+00	4.935543e+02
3.480000e+02	4.943947e+02	4.319771e+02	2.081476e+01	3.623896e+01	1.442776e+00	7.540347e-02	3.845680e+00	0.000000e+00	4.943947e+02
3.490000e+02	5.006141e+02	4.387307e+02	2.136945e+01	3.537660e+01	1.391786e+00	7.775486e-02	3.667792e+00	0.000000e+00	5.006141e+02
3.500000e+02	5.029466e+02	4.454815e+02	1.543572e+01	3.698864e+01	1.327284e+00	8.010625e-02	3.633370e+00	0.000000e+00	5.029466e+02
3.510000e+02	4.998736e+02	4.411576e+02	1.549612e+01	3.825853e+01	1.270779e+00	8.150942e-02	3.609096e+00	0.000000e+00	4.998736e+02
3.520000e+02	4.817221e+02	4.201552e+02	1.601390e+01	4.067367e+01	1.214275e+00	8.410277e-02	3.580939e+00	0.000000e+00	4.817221e+02
3.530000e+02	4.760784e+02	4.125679e+02	1.652242e+01	4.218435e+01	1.165140e+00	8.436287e-02	3.554284e+00	0.000000e+00	4.760784e+02
3.540000e+02	4.615007e+02	3.967289e+02	1.669197e+01	4.353408e+01	1.085297e+00	8.697044e-02	3.373484e+00	0.000000e+00	4.615007e+02
3.550000e+02	4.657009e+02	4.013952e+02	1.726802e+01	4.273754e+01	1.021422e+00	8.843492e-02	3.190303e+00	0.000000e+00	4.657009e+02
3.560000e+02	4.713097e+02	4.047459e+02	1.783238e+01	4.449235e+01	9.808860e-01	8.868241e-02	3.169474e+00	0.000000e+00	4.713097e+02
3.570000e+02	4.322859e+02	3.662397e+02	1.780710e+01	4.421277e+01	9.397226e-01	9.006582e-02	2.996534e+00	0.000000e+00	4.322859e+02
3.580000e+02	4.485332e+02	3.725479e+02	1.799542e+01	4.651638e+01	5.828599e+00	8.506544e-02	5.559828e+00	0.000000e+00	4.485332e+02
3.590000e+02	4.438977e+02	3.779038e+02	1.679298e+01	4.469647e+01	1.270625e+00	8.388975e-02	3.149943e+00	0.000000e+00	4.438977e+02
3.600000e+02	4.525286e+02	3.842864e+02	1.706239e+01	4.659812e+01	1.289867e+00	8.741683e-02	3.204373e+00	0.000000e+00	4.525286e+02
3.610000e+02	4.582440e+02	3.872516e+02	1.755142e+01	4.898193e+01	1.320156e+00	8.741683e-02	3.051466e+00	0.000000e+00	4.582440e+02
3.620000e+02	4.663131e+02	3.938127e+02	1.818505e+01	4.975003e+01	1.311268e+00	9.094391e-02	3.163052e+00	0.000000e+00	4.663131e+02
3.630000e+02	4.652810e+02	3.941207e+02	1.857253e+01	4.800406e+01	1.305168e+00	8.859252e-02	3.189878e+00	0.000000e+00	4.652810e+02
3.640000e+02	4.624339e+02	3.919782e+02	1.862329e+01	4.661051e+01	1.269471e+00	9.101678e-02	3.861433e+00	0.000000e+00	4.624339e+02
3.650000e+02	4.673216e+02	3.981866e+02	1.915330e+01	4.401069e+01	1.124060e+00	9.101678e-02	4.755932e+00	0.000000e+00	4.673216e+02
3.660000e+02	4.757858e+02	4.047006e+02	1.990632e+01	4.427790e+01	9.869294e-01	9.094391e-02	5.823059e+00	0.000000e+00	4.757858e+02
3.670000e+02	4.829437e+02	4.099253e+02	2.061586e+01	4.434171e+01	8.959578e-01	8.976822e-02	7.075071e+00	0.000000e+00	4.829437e+02
3.680000e+02	4.923823e+02	4.164911e+02	1.985805e+01	4.632722e+01	8.677055e-01	8.859252e-02	8.749611e+00	0.000000e+00	4.923823e+02
3.690000e+02	4.850531e+02	4.093103e+02	2.051775e+01	4.684610e+01	8.405632e-01	8.976822e-02	7.448598e+00	0.000000e+00	4.850531e+02
3.700000e+02	4.745518e+02	4.019127e+02	2.075470e+01	4.465035e+01	7.770069e-01	8.859252e-02	6.368392e+00	0.000000e+00	4.745518e+02
3.710000e+02	4.663131e+02	3.890591e+02	2.103757e+01	4.654056e+01	2.775432e+00	8.741683e-02	6.812950e+00	0.000000e+00	4.663131e+02
3.720000e+02	4.712093e+02	3.958357e+02	2.077851e+01	4.747335e+01	1.096817e+00	8.388975e-02	5.941042e+00	0.000000e+00	4.712093e+02
3.730000e+02	4.787235e+02	4.028047e+02	2.107259e+01	4.825484e+01	1.049348e+00	8.506544e-02	5.456953e+00	0.000000e+00	4.787235e+02
3.740000e+02	4.854174e+02	4.094552e+02	2.173904e+01	4.785359e+01	9.950636e-01	8.741683e-02	5.287175e+00	0.000000e+00	4.854174e+02
3.750000e+02	4.929227e+02	4.159753e+02	2.246327e+01	4.848816e+01	9.473576e-01	8.741683e-02	4.961212e+00	0.000000e+00	4.929227e+02
3.760000e+02	4.665603e+02	3.874076e+02	2.314144e+01	5.007743e+01	9.048017e-01	8.859252e-02	4.940384e+00	0.000000e+00	4.665603e+02
3.770000e+02	4.751537e+02	3.942697e+02	2.391694e+01	5.108599e+01	8.614542e-01	9.094391e-02	4.928732e+00	0.000000e+00	4.751537e+02
3.780000e+02	4.524420e+02	3.728193e+02	2.246242e+01	5.134994e+01	8.077247e-01	9.329530e-02	4.909313e+00	0.000000e+00	4.524420e+02
3.790000e+02	4.573689e+02	3.784080e+02	2.327907e+01	5.007518e+01	7.732123e-01	9.094391e-02	4.742448e+00	0.000000e+00	4.573689e+02
3.800000e+02	4.642589e+02	3.856501e+02	2.410352e+01	4.908919e+01	7.492001e-01	8.976822e-02	4.577183e+00	0.000000e+00	4.642589e+02
3.810000e+02	4.510061e+02	3.729460e+02	2.471509e+01	4.796892e+01	7.208295e-01	8.976822e-02	4.565532e+00	0.000000e+00	4.510061e+02
3.820000e+02	4.549354e+02	3.759835e+02	2.554953e+01	4.806441e+01	6.912305e-01	9.094391e-02	4.555822e+00	0.000000e+00	4.549354e+02
3.830000e+02	4.569288e+02	3.775246e+02	2.633167e+01	4.824186e+01	6.571549e-01	9.211961e-02	4.081443e+00	0.000000e+00	4.569288e+02
3.840000e+02	4.642467e+02	3.845261e+02	2.543694e+01	4.950281e+01	6.158273e-01	9.329530e-02	4.071733e+00	0.000000e+00	4.642467e+02
3.850000e+02	4.712711e+02	3.920315e+02	2.624723e+01	4.876774e+01	5.499325e-01	9.474396e-02	3.579877e+00	0.000000e+00	4.712711e+02
3.860000e+02	4.758479e+02	3.973072e+02	2.723347e+01	4.693254e+01	7.463520e-01	9.620083e-02	3.532096e+00	0.000000e+00	4.758479e+02
3.870000e+02	4.732200e+02	3.965959e+02	2.790624e+01	4.459212e+01	6.848156e-01	9.414501e-02	3.346783e+00	0.000000e+00	4.732200e+02
3.880000e+02	4.766813e+02	4.007554e+02	2.748852e+01	4.450726e+01	6.576734e-01	9.447100e-02	3.177976e+00	0.000000e+00	4.766813e+02
3.890000e+02	4.842323e+02	4.076439e+02	2.757031e+01	4.559164e+01	6.286294e-01	9.329530e-02	2.704567e+00	0.000000e+00	4.842323e+02
3.900000e+02	4.606518e+02	3.871719e+02	2.758411e+01	4.267460e+01	5.954637e-01	9.094391e-02	2.534789e+00	0.000000e+00	4.606518e+02
3.910000e+02	4.636093e+02	3.903333e+02	2.707748e+01	4.322841e+01	5.296872e-01	9.094391e-02	2.349476e+00	0.000000e+00	4.636093e+02
3.920000e+02	4.731167e+02	3.982745e+02	2.793164e+01	4.411761e+01	5.088051e-01	9.211961e-02	2.191979e+00	0.000000e+00	4.731167e+02
3.930000e+02	4.829680e+02	4.063074e+02	2.881895e+01	4.508916e+01	4.842379e-01	8.506544e-02	2.183240e+00	0.000000e+00	4.829680e+02
3.940000e+02	4.858999e+02	4.091144e+02	2.980218e+01	4.425875e+01	4.645841e-01	8.741683e-02	2.172560e+00	0.000000e+00	4.858999e+02
3.950000e+02	4.873320e+02	4.122205e+02	3.082703e+01	4.174442e+01	4.437020e-01	8.388975e-02	2.012491e+00	0.000000e+00	4.873320e+02
3.960000e+02	4.969574e+02	4.198608e+02	3.188377e+01	4.269434e+01	4.270600e-01	8.859252e-02	2.002782e+00	0.000000e+00	4.969574e+02
3.970000e+02	5.001694e+02	4.247063e+02	3.218234e+01	4.079258e+01	4.067329e-01	8.741683e-02	1.994043e+00	0.000000e+00	5.001694e+02
3.980000e+02	4.905805e+02	4.152978e+02	3.160375e+01	4.151285e+01	3.937759e-01	9.094391e-02	1.681332e+00	0.000000e+00	4.905805e+02
3.990000e+02	4.923547e+02	4.178032e+02	3.084333e+01	3.863625e+01	2.299400e+00	8.624114e-02	2.686260e+00	0.000000e+00	4.923547e+02
4.000000e+02	4.994430e+02	4.261204e+02	3.170556e+01	3.894517e+01	7.209566e-01	8.506544e-02	1.865812e+00	0.000000e+00	4.994430e+02
